LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY ALU2 IS
PORT(
	Clock : IN STD_LOGIC; -- input clock signal
	A,B : IN UNSIGNED(7 DOWNTO 0); -- 8 bit inputs from latches A and B
	student_id : IN UNSIGNED (3 DOWNTO 0); --4 bit student id from FSM
	OP : IN UNSIGNED(15 DOWNTO 0); -- 16 bit selector for Operation from Decoder
	Neg : OUT STD_LOGIC; -- is the result negative? set-ve bit output
	R1 : OUT UNSIGNED (3 DOWNTO 0); -- lower 4 bits of 8 bit Result Output 
	R2 : OUT UNSIGNED (3 DOWNTO 0)); -- higher 4 bits of 8-bit Result Output 
END ALU2;

ARCHITECTURE calculation OF ALU2 IS
SIGNAL Reg1, Reg2, Result : UNSIGNED(7 DOWNTO 0):= (OTHERS =>'0');
SIGNAL Reg4 : UNSIGNED(0 TO 7);
SIGNAL temp : STD_LOGIC;
BEGIN 
Reg1 <= A; -- temporarily stores A in Reg1 local variable 
Reg2 <= B; -- temporarily stores B in Reg2 local variable 
PROCESS(Clock, OP)
BEGIN 
	IF(rising_edge(Clock)) THEN --Do the calculation @ positive edge of clock cycle 
		CASE OP IS
			WHEN "0000000000000001"=> -- Difference Between A and B
				Result <= Reg1 + (not(Reg2)+1);
				Neg <= '0';
			WHEN "0000000000000010"=> -- 2's Complement of B
				Result <= (not(Reg2)+1);
				Neg <= '0';
			WHEN "0000000000000100"=> -- Swap lower bits of A with lower bits of B
				Result <= Reg1(7 DOWNTO 4) & Reg2(3 DOWNTO 0);
				Neg <= '0';
			WHEN "0000000000001000"=> -- Null on output
				Result <= null;
				Neg <= null;
			WHEN "0000000000010000"=> -- Decrement B by 5
				Result <= (Reg2 - 5);
				Neg <= '0';
			WHEN "0000000000100000"=> -- Invert bit-significance order of A 
				Result <= Reg1;
				Neg<= '1';
			WHEN "0000000001000000"=>-- Shift B to left by 3 bits, input bit = 1 (SHL) 
				--temp <= Reg2(7);
				Result(7) <= Reg2(6);
				Result(6) <= Reg2(5);
				Result(5) <= Reg2(4);
				Result(4) <= Reg2(3);
				Result(3) <= Reg2(2);
				Result(2) <= Reg2(1);
				Result(1) <= Reg2(0);
				Result(0) <= '1';
				Neg <= '0';
			WHEN "0000000010000000"=> -- Increment A by 3
				Result <= (Reg1 + 3);
				Neg <= '0';
			WHEN "0000000100000000"=> -- Invert All Bits of B
				Result(7) <= Reg2(0);
				Result(6) <= Reg2(1);
				Result(5) <= Reg2(2);
				Result(4) <= Reg2(3);
				Result(3) <= Reg2(4);
				Result(2) <= Reg2(5);
				Result(1) <= Reg2(6);
				Result(0) <= Reg2(7);
				Neg <= '0';
			WHEN OTHERS =>
				Result <= "00000000";
				Neg <= '0';
		END CASE;
	END IF;
END PROCESS;
R1 <= Result(3 DOWNTO 0);
R2 <= Result(7 DOWNTO 4);
END calculation;